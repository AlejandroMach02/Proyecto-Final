----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 17.03.2024 13:12:00
-- Design Name: 
-- Module Name: conta_generic - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity conta_generic is
  generic ( 
    fin_conta: natural := 10**7;                -- frecuencia inicial es 100MHz y queremos la f de 1 decima de segundo, la nueva frecuencia ser� de 10*10e6
    n_bits: natural := 24;                      -- la menos potencia de 2 superior a 10e6 es 24 -->2^3<10e6<2^4
    max: unsigned:="1001");
  Port ( 
    clk: in std_logic;
    rst: in std_logic;
    enable: in std_logic;                       -- se�al del contador anterior
    up_down: in std_logic;                      -- interruptor de cuenta ascendente/descendente SW OFF = ASCENDENTE, SW ON= DESCENDENTE
    sconta: out std_logic;                      -- emitir� una se�al/pulso cada periodo, si es s1dec, emirtira un pulso cada decima de segundo, si es s1seg emitira un un pulso cada segundo.. 
    vconta: out unsigned (n_bits-1 downto 0));  -- tendr� los bits necesarios para contar hasta el valor deseado y mostrarlo luego en los displays. se realiza a partir de la se�al s-conta. 
end conta_generic;

architecture Behavioral of conta_generic is

-- se�ales intermedias
    signal contador: unsigned (n_bits-1 downto 0);  -- se�al que lleva la cuenta, debe tener un rango potencia de 2. 
    signal s_conta : std_logic;
   
begin

P_contageneric: process (clk, rst)       -- descripcion del contador
begin
    if rst ='1' then
        contador <= (others=>'0');
    elsif clk'event and clk='1' then
        if enable='1' then 
            if up_down ='0' then   
                if s_conta='1' then
                contador<=(others=>'0');
                else
                contador<=contador + 1;
                end if;
            else   -- si up_down esta en 1 
                if s_conta='1' then
                contador<=max;
                else
                contador<=contador-1;
                end if;
            end if;
        end if;
    end if;
end process;

s_conta<= '1' when contador = fin_conta-1 and enable ='1' and up_down='0' else
          '1' when contador = 0 and enable ='1' and up_down ='1' else '0';  
sconta<=s_conta;
vconta<=contador;

end Behavioral;